// nios_flash_interface.v

// Generated using ACDS version 13.0sp1 232 at 2018.02.05.15:56:54

`timescale 1 ps / 1 ps
module nios_flash_interface (
		input  wire  clock_50_clk,               //              clock_50.clk
		input  wire  reset_n_reset_n,            //               reset_n.reset_n
		input  wire  spi_mediator_external_MISO, // spi_mediator_external.MISO
		output wire  spi_mediator_external_MOSI, //                      .MOSI
		output wire  spi_mediator_external_SCLK, //                      .SCLK
		output wire  spi_mediator_external_SS_n  //                      .SS_n
	);

	wire         niosii_instruction_master_waitrequest;                                                              // NIOSII_instruction_master_translator:av_waitrequest -> NIOSII:i_waitrequest
	wire  [25:0] niosii_instruction_master_address;                                                                  // NIOSII:i_address -> NIOSII_instruction_master_translator:av_address
	wire         niosii_instruction_master_read;                                                                     // NIOSII:i_read -> NIOSII_instruction_master_translator:av_read
	wire  [31:0] niosii_instruction_master_readdata;                                                                 // NIOSII_instruction_master_translator:av_readdata -> NIOSII:i_readdata
	wire         niosii_data_master_waitrequest;                                                                     // NIOSII_data_master_translator:av_waitrequest -> NIOSII:d_waitrequest
	wire  [31:0] niosii_data_master_writedata;                                                                       // NIOSII:d_writedata -> NIOSII_data_master_translator:av_writedata
	wire  [25:0] niosii_data_master_address;                                                                         // NIOSII:d_address -> NIOSII_data_master_translator:av_address
	wire         niosii_data_master_write;                                                                           // NIOSII:d_write -> NIOSII_data_master_translator:av_write
	wire         niosii_data_master_read;                                                                            // NIOSII:d_read -> NIOSII_data_master_translator:av_read
	wire  [31:0] niosii_data_master_readdata;                                                                        // NIOSII_data_master_translator:av_readdata -> NIOSII:d_readdata
	wire         niosii_data_master_debugaccess;                                                                     // NIOSII:jtag_debug_module_debugaccess_to_roms -> NIOSII_data_master_translator:av_debugaccess
	wire   [3:0] niosii_data_master_byteenable;                                                                      // NIOSII:d_byteenable -> NIOSII_data_master_translator:av_byteenable
	wire         niosii_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest;                                // NIOSII:jtag_debug_module_waitrequest -> NIOSII_jtag_debug_module_translator:av_waitrequest
	wire  [31:0] niosii_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                  // NIOSII_jtag_debug_module_translator:av_writedata -> NIOSII:jtag_debug_module_writedata
	wire   [8:0] niosii_jtag_debug_module_translator_avalon_anti_slave_0_address;                                    // NIOSII_jtag_debug_module_translator:av_address -> NIOSII:jtag_debug_module_address
	wire         niosii_jtag_debug_module_translator_avalon_anti_slave_0_write;                                      // NIOSII_jtag_debug_module_translator:av_write -> NIOSII:jtag_debug_module_write
	wire         niosii_jtag_debug_module_translator_avalon_anti_slave_0_read;                                       // NIOSII_jtag_debug_module_translator:av_read -> NIOSII:jtag_debug_module_read
	wire  [31:0] niosii_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                   // NIOSII:jtag_debug_module_readdata -> NIOSII_jtag_debug_module_translator:av_readdata
	wire         niosii_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                // NIOSII_jtag_debug_module_translator:av_debugaccess -> NIOSII:jtag_debug_module_debugaccess
	wire   [3:0] niosii_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                 // NIOSII_jtag_debug_module_translator:av_byteenable -> NIOSII:jtag_debug_module_byteenable
	wire         bridge_s0_translator_avalon_anti_slave_0_waitrequest;                                               // BRIDGE:s0_waitrequest -> BRIDGE_s0_translator:av_waitrequest
	wire   [0:0] bridge_s0_translator_avalon_anti_slave_0_burstcount;                                                // BRIDGE_s0_translator:av_burstcount -> BRIDGE:s0_burstcount
	wire  [31:0] bridge_s0_translator_avalon_anti_slave_0_writedata;                                                 // BRIDGE_s0_translator:av_writedata -> BRIDGE:s0_writedata
	wire  [15:0] bridge_s0_translator_avalon_anti_slave_0_address;                                                   // BRIDGE_s0_translator:av_address -> BRIDGE:s0_address
	wire         bridge_s0_translator_avalon_anti_slave_0_write;                                                     // BRIDGE_s0_translator:av_write -> BRIDGE:s0_write
	wire         bridge_s0_translator_avalon_anti_slave_0_read;                                                      // BRIDGE_s0_translator:av_read -> BRIDGE:s0_read
	wire  [31:0] bridge_s0_translator_avalon_anti_slave_0_readdata;                                                  // BRIDGE:s0_readdata -> BRIDGE_s0_translator:av_readdata
	wire         bridge_s0_translator_avalon_anti_slave_0_debugaccess;                                               // BRIDGE_s0_translator:av_debugaccess -> BRIDGE:s0_debugaccess
	wire         bridge_s0_translator_avalon_anti_slave_0_readdatavalid;                                             // BRIDGE:s0_readdatavalid -> BRIDGE_s0_translator:av_readdatavalid
	wire   [3:0] bridge_s0_translator_avalon_anti_slave_0_byteenable;                                                // BRIDGE_s0_translator:av_byteenable -> BRIDGE:s0_byteenable
	wire   [0:0] bridge_m0_burstcount;                                                                               // BRIDGE:m0_burstcount -> BRIDGE_m0_translator:av_burstcount
	wire         bridge_m0_waitrequest;                                                                              // BRIDGE_m0_translator:av_waitrequest -> BRIDGE:m0_waitrequest
	wire  [15:0] bridge_m0_address;                                                                                  // BRIDGE:m0_address -> BRIDGE_m0_translator:av_address
	wire  [31:0] bridge_m0_writedata;                                                                                // BRIDGE:m0_writedata -> BRIDGE_m0_translator:av_writedata
	wire         bridge_m0_write;                                                                                    // BRIDGE:m0_write -> BRIDGE_m0_translator:av_write
	wire         bridge_m0_read;                                                                                     // BRIDGE:m0_read -> BRIDGE_m0_translator:av_read
	wire  [31:0] bridge_m0_readdata;                                                                                 // BRIDGE_m0_translator:av_readdata -> BRIDGE:m0_readdata
	wire         bridge_m0_debugaccess;                                                                              // BRIDGE:m0_debugaccess -> BRIDGE_m0_translator:av_debugaccess
	wire   [3:0] bridge_m0_byteenable;                                                                               // BRIDGE:m0_byteenable -> BRIDGE_m0_translator:av_byteenable
	wire         bridge_m0_readdatavalid;                                                                            // BRIDGE_m0_translator:av_readdatavalid -> BRIDGE:m0_readdatavalid
	wire  [31:0] onchip_ram_s1_translator_avalon_anti_slave_0_writedata;                                             // ONCHIP_RAM_s1_translator:av_writedata -> ONCHIP_RAM:writedata
	wire   [9:0] onchip_ram_s1_translator_avalon_anti_slave_0_address;                                               // ONCHIP_RAM_s1_translator:av_address -> ONCHIP_RAM:address
	wire         onchip_ram_s1_translator_avalon_anti_slave_0_chipselect;                                            // ONCHIP_RAM_s1_translator:av_chipselect -> ONCHIP_RAM:chipselect
	wire         onchip_ram_s1_translator_avalon_anti_slave_0_clken;                                                 // ONCHIP_RAM_s1_translator:av_clken -> ONCHIP_RAM:clken
	wire         onchip_ram_s1_translator_avalon_anti_slave_0_write;                                                 // ONCHIP_RAM_s1_translator:av_write -> ONCHIP_RAM:write
	wire  [31:0] onchip_ram_s1_translator_avalon_anti_slave_0_readdata;                                              // ONCHIP_RAM:readdata -> ONCHIP_RAM_s1_translator:av_readdata
	wire   [3:0] onchip_ram_s1_translator_avalon_anti_slave_0_byteenable;                                            // ONCHIP_RAM_s1_translator:av_byteenable -> ONCHIP_RAM:byteenable
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                             // JTAG_UART:av_waitrequest -> JTAG_UART_avalon_jtag_slave_translator:av_waitrequest
	wire  [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                               // JTAG_UART_avalon_jtag_slave_translator:av_writedata -> JTAG_UART:av_writedata
	wire   [0:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                 // JTAG_UART_avalon_jtag_slave_translator:av_address -> JTAG_UART:av_address
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                              // JTAG_UART_avalon_jtag_slave_translator:av_chipselect -> JTAG_UART:av_chipselect
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                   // JTAG_UART_avalon_jtag_slave_translator:av_write -> JTAG_UART:av_write_n
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                    // JTAG_UART_avalon_jtag_slave_translator:av_read -> JTAG_UART:av_read_n
	wire  [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                // JTAG_UART:av_readdata -> JTAG_UART_avalon_jtag_slave_translator:av_readdata
	wire  [15:0] timer_s1_translator_avalon_anti_slave_0_writedata;                                                  // TIMER_s1_translator:av_writedata -> TIMER:writedata
	wire   [2:0] timer_s1_translator_avalon_anti_slave_0_address;                                                    // TIMER_s1_translator:av_address -> TIMER:address
	wire         timer_s1_translator_avalon_anti_slave_0_chipselect;                                                 // TIMER_s1_translator:av_chipselect -> TIMER:chipselect
	wire         timer_s1_translator_avalon_anti_slave_0_write;                                                      // TIMER_s1_translator:av_write -> TIMER:write_n
	wire  [15:0] timer_s1_translator_avalon_anti_slave_0_readdata;                                                   // TIMER:readdata -> TIMER_s1_translator:av_readdata
	wire  [15:0] spi_mediator_spi_control_port_translator_avalon_anti_slave_0_writedata;                             // SPI_MEDIATOR_spi_control_port_translator:av_writedata -> SPI_MEDIATOR:data_from_cpu
	wire   [2:0] spi_mediator_spi_control_port_translator_avalon_anti_slave_0_address;                               // SPI_MEDIATOR_spi_control_port_translator:av_address -> SPI_MEDIATOR:mem_addr
	wire         spi_mediator_spi_control_port_translator_avalon_anti_slave_0_chipselect;                            // SPI_MEDIATOR_spi_control_port_translator:av_chipselect -> SPI_MEDIATOR:spi_select
	wire         spi_mediator_spi_control_port_translator_avalon_anti_slave_0_write;                                 // SPI_MEDIATOR_spi_control_port_translator:av_write -> SPI_MEDIATOR:write_n
	wire         spi_mediator_spi_control_port_translator_avalon_anti_slave_0_read;                                  // SPI_MEDIATOR_spi_control_port_translator:av_read -> SPI_MEDIATOR:read_n
	wire  [15:0] spi_mediator_spi_control_port_translator_avalon_anti_slave_0_readdata;                              // SPI_MEDIATOR:data_to_cpu -> SPI_MEDIATOR_spi_control_port_translator:av_readdata
	wire         niosii_instruction_master_translator_avalon_universal_master_0_waitrequest;                         // NIOSII_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> NIOSII_instruction_master_translator:uav_waitrequest
	wire   [2:0] niosii_instruction_master_translator_avalon_universal_master_0_burstcount;                          // NIOSII_instruction_master_translator:uav_burstcount -> NIOSII_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] niosii_instruction_master_translator_avalon_universal_master_0_writedata;                           // NIOSII_instruction_master_translator:uav_writedata -> NIOSII_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [25:0] niosii_instruction_master_translator_avalon_universal_master_0_address;                             // NIOSII_instruction_master_translator:uav_address -> NIOSII_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         niosii_instruction_master_translator_avalon_universal_master_0_lock;                                // NIOSII_instruction_master_translator:uav_lock -> NIOSII_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         niosii_instruction_master_translator_avalon_universal_master_0_write;                               // NIOSII_instruction_master_translator:uav_write -> NIOSII_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         niosii_instruction_master_translator_avalon_universal_master_0_read;                                // NIOSII_instruction_master_translator:uav_read -> NIOSII_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] niosii_instruction_master_translator_avalon_universal_master_0_readdata;                            // NIOSII_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> NIOSII_instruction_master_translator:uav_readdata
	wire         niosii_instruction_master_translator_avalon_universal_master_0_debugaccess;                         // NIOSII_instruction_master_translator:uav_debugaccess -> NIOSII_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] niosii_instruction_master_translator_avalon_universal_master_0_byteenable;                          // NIOSII_instruction_master_translator:uav_byteenable -> NIOSII_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         niosii_instruction_master_translator_avalon_universal_master_0_readdatavalid;                       // NIOSII_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> NIOSII_instruction_master_translator:uav_readdatavalid
	wire         niosii_data_master_translator_avalon_universal_master_0_waitrequest;                                // NIOSII_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> NIOSII_data_master_translator:uav_waitrequest
	wire   [2:0] niosii_data_master_translator_avalon_universal_master_0_burstcount;                                 // NIOSII_data_master_translator:uav_burstcount -> NIOSII_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] niosii_data_master_translator_avalon_universal_master_0_writedata;                                  // NIOSII_data_master_translator:uav_writedata -> NIOSII_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [25:0] niosii_data_master_translator_avalon_universal_master_0_address;                                    // NIOSII_data_master_translator:uav_address -> NIOSII_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         niosii_data_master_translator_avalon_universal_master_0_lock;                                       // NIOSII_data_master_translator:uav_lock -> NIOSII_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         niosii_data_master_translator_avalon_universal_master_0_write;                                      // NIOSII_data_master_translator:uav_write -> NIOSII_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         niosii_data_master_translator_avalon_universal_master_0_read;                                       // NIOSII_data_master_translator:uav_read -> NIOSII_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] niosii_data_master_translator_avalon_universal_master_0_readdata;                                   // NIOSII_data_master_translator_avalon_universal_master_0_agent:av_readdata -> NIOSII_data_master_translator:uav_readdata
	wire         niosii_data_master_translator_avalon_universal_master_0_debugaccess;                                // NIOSII_data_master_translator:uav_debugaccess -> NIOSII_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] niosii_data_master_translator_avalon_universal_master_0_byteenable;                                 // NIOSII_data_master_translator:uav_byteenable -> NIOSII_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         niosii_data_master_translator_avalon_universal_master_0_readdatavalid;                              // NIOSII_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> NIOSII_data_master_translator:uav_readdatavalid
	wire         niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                  // NIOSII_jtag_debug_module_translator:uav_waitrequest -> NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                   // NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> NIOSII_jtag_debug_module_translator:uav_burstcount
	wire  [31:0] niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                    // NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> NIOSII_jtag_debug_module_translator:uav_writedata
	wire  [25:0] niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                      // NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> NIOSII_jtag_debug_module_translator:uav_address
	wire         niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                        // NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> NIOSII_jtag_debug_module_translator:uav_write
	wire         niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                         // NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> NIOSII_jtag_debug_module_translator:uav_lock
	wire         niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                         // NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> NIOSII_jtag_debug_module_translator:uav_read
	wire  [31:0] niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                     // NIOSII_jtag_debug_module_translator:uav_readdata -> NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                // NIOSII_jtag_debug_module_translator:uav_readdatavalid -> NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                  // NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> NIOSII_jtag_debug_module_translator:uav_debugaccess
	wire   [3:0] niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                   // NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> NIOSII_jtag_debug_module_translator:uav_byteenable
	wire         niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;           // NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                 // NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;         // NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                  // NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                 // NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;        // NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;              // NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;      // NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;               // NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;              // NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;            // NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;             // NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;            // NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // BRIDGE_s0_translator:uav_waitrequest -> BRIDGE_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // BRIDGE_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> BRIDGE_s0_translator:uav_burstcount
	wire  [31:0] bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // BRIDGE_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> BRIDGE_s0_translator:uav_writedata
	wire  [25:0] bridge_s0_translator_avalon_universal_slave_0_agent_m0_address;                                     // BRIDGE_s0_translator_avalon_universal_slave_0_agent:m0_address -> BRIDGE_s0_translator:uav_address
	wire         bridge_s0_translator_avalon_universal_slave_0_agent_m0_write;                                       // BRIDGE_s0_translator_avalon_universal_slave_0_agent:m0_write -> BRIDGE_s0_translator:uav_write
	wire         bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock;                                        // BRIDGE_s0_translator_avalon_universal_slave_0_agent:m0_lock -> BRIDGE_s0_translator:uav_lock
	wire         bridge_s0_translator_avalon_universal_slave_0_agent_m0_read;                                        // BRIDGE_s0_translator_avalon_universal_slave_0_agent:m0_read -> BRIDGE_s0_translator:uav_read
	wire  [31:0] bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // BRIDGE_s0_translator:uav_readdata -> BRIDGE_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // BRIDGE_s0_translator:uav_readdatavalid -> BRIDGE_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // BRIDGE_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> BRIDGE_s0_translator:uav_debugaccess
	wire   [3:0] bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // BRIDGE_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> BRIDGE_s0_translator:uav_byteenable
	wire         bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // BRIDGE_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> BRIDGE_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // BRIDGE_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> BRIDGE_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // BRIDGE_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> BRIDGE_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [95:0] bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // BRIDGE_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> BRIDGE_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // BRIDGE_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> BRIDGE_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // BRIDGE_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> BRIDGE_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // BRIDGE_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> BRIDGE_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // BRIDGE_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> BRIDGE_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [95:0] bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // BRIDGE_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> BRIDGE_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // BRIDGE_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> BRIDGE_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // BRIDGE_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> BRIDGE_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // BRIDGE_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> BRIDGE_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // BRIDGE_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> BRIDGE_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         bridge_m0_translator_avalon_universal_master_0_waitrequest;                                         // BRIDGE_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> BRIDGE_m0_translator:uav_waitrequest
	wire   [2:0] bridge_m0_translator_avalon_universal_master_0_burstcount;                                          // BRIDGE_m0_translator:uav_burstcount -> BRIDGE_m0_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] bridge_m0_translator_avalon_universal_master_0_writedata;                                           // BRIDGE_m0_translator:uav_writedata -> BRIDGE_m0_translator_avalon_universal_master_0_agent:av_writedata
	wire  [15:0] bridge_m0_translator_avalon_universal_master_0_address;                                             // BRIDGE_m0_translator:uav_address -> BRIDGE_m0_translator_avalon_universal_master_0_agent:av_address
	wire         bridge_m0_translator_avalon_universal_master_0_lock;                                                // BRIDGE_m0_translator:uav_lock -> BRIDGE_m0_translator_avalon_universal_master_0_agent:av_lock
	wire         bridge_m0_translator_avalon_universal_master_0_write;                                               // BRIDGE_m0_translator:uav_write -> BRIDGE_m0_translator_avalon_universal_master_0_agent:av_write
	wire         bridge_m0_translator_avalon_universal_master_0_read;                                                // BRIDGE_m0_translator:uav_read -> BRIDGE_m0_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] bridge_m0_translator_avalon_universal_master_0_readdata;                                            // BRIDGE_m0_translator_avalon_universal_master_0_agent:av_readdata -> BRIDGE_m0_translator:uav_readdata
	wire         bridge_m0_translator_avalon_universal_master_0_debugaccess;                                         // BRIDGE_m0_translator:uav_debugaccess -> BRIDGE_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] bridge_m0_translator_avalon_universal_master_0_byteenable;                                          // BRIDGE_m0_translator:uav_byteenable -> BRIDGE_m0_translator_avalon_universal_master_0_agent:av_byteenable
	wire         bridge_m0_translator_avalon_universal_master_0_readdatavalid;                                       // BRIDGE_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> BRIDGE_m0_translator:uav_readdatavalid
	wire         onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // ONCHIP_RAM_s1_translator:uav_waitrequest -> ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ONCHIP_RAM_s1_translator:uav_burstcount
	wire  [31:0] onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                               // ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ONCHIP_RAM_s1_translator:uav_writedata
	wire  [15:0] onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_address;                                 // ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:m0_address -> ONCHIP_RAM_s1_translator:uav_address
	wire         onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_write;                                   // ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:m0_write -> ONCHIP_RAM_s1_translator:uav_write
	wire         onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                    // ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ONCHIP_RAM_s1_translator:uav_lock
	wire         onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_read;                                    // ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:m0_read -> ONCHIP_RAM_s1_translator:uav_read
	wire  [31:0] onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                // ONCHIP_RAM_s1_translator:uav_readdata -> ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // ONCHIP_RAM_s1_translator:uav_readdatavalid -> ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ONCHIP_RAM_s1_translator:uav_debugaccess
	wire   [3:0] onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ONCHIP_RAM_s1_translator:uav_byteenable
	wire         onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [85:0] onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                             // ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [85:0] onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         onchip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] onchip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         onchip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;               // JTAG_UART_avalon_jtag_slave_translator:uav_waitrequest -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> JTAG_UART_avalon_jtag_slave_translator:uav_burstcount
	wire  [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                 // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> JTAG_UART_avalon_jtag_slave_translator:uav_writedata
	wire  [15:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                   // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> JTAG_UART_avalon_jtag_slave_translator:uav_address
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                     // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> JTAG_UART_avalon_jtag_slave_translator:uav_write
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                      // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> JTAG_UART_avalon_jtag_slave_translator:uav_lock
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                      // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> JTAG_UART_avalon_jtag_slave_translator:uav_read
	wire  [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                  // JTAG_UART_avalon_jtag_slave_translator:uav_readdata -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;             // JTAG_UART_avalon_jtag_slave_translator:uav_readdatavalid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;               // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> JTAG_UART_avalon_jtag_slave_translator:uav_debugaccess
	wire   [3:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> JTAG_UART_avalon_jtag_slave_translator:uav_byteenable
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;        // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;              // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;      // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [85:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;               // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;              // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;     // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;           // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;   // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [85:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;            // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;           // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;         // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;          // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;         // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // TIMER_s1_translator:uav_waitrequest -> TIMER_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // TIMER_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> TIMER_s1_translator:uav_burstcount
	wire  [31:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // TIMER_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> TIMER_s1_translator:uav_writedata
	wire  [15:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // TIMER_s1_translator_avalon_universal_slave_0_agent:m0_address -> TIMER_s1_translator:uav_address
	wire         timer_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // TIMER_s1_translator_avalon_universal_slave_0_agent:m0_write -> TIMER_s1_translator:uav_write
	wire         timer_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // TIMER_s1_translator_avalon_universal_slave_0_agent:m0_lock -> TIMER_s1_translator:uav_lock
	wire         timer_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // TIMER_s1_translator_avalon_universal_slave_0_agent:m0_read -> TIMER_s1_translator:uav_read
	wire  [31:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // TIMER_s1_translator:uav_readdata -> TIMER_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // TIMER_s1_translator:uav_readdatavalid -> TIMER_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // TIMER_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> TIMER_s1_translator:uav_debugaccess
	wire   [3:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // TIMER_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> TIMER_s1_translator:uav_byteenable
	wire         timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // TIMER_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> TIMER_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // TIMER_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> TIMER_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // TIMER_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> TIMER_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [85:0] timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // TIMER_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> TIMER_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // TIMER_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> TIMER_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // TIMER_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> TIMER_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // TIMER_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> TIMER_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // TIMER_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> TIMER_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [85:0] timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // TIMER_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> TIMER_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // TIMER_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> TIMER_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // TIMER_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> TIMER_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // TIMER_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> TIMER_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // TIMER_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> TIMER_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // SPI_MEDIATOR_spi_control_port_translator:uav_waitrequest -> SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount;              // SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:m0_burstcount -> SPI_MEDIATOR_spi_control_port_translator:uav_burstcount
	wire  [31:0] spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata;               // SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:m0_writedata -> SPI_MEDIATOR_spi_control_port_translator:uav_writedata
	wire  [15:0] spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address;                 // SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:m0_address -> SPI_MEDIATOR_spi_control_port_translator:uav_address
	wire         spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write;                   // SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:m0_write -> SPI_MEDIATOR_spi_control_port_translator:uav_write
	wire         spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock;                    // SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:m0_lock -> SPI_MEDIATOR_spi_control_port_translator:uav_lock
	wire         spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read;                    // SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:m0_read -> SPI_MEDIATOR_spi_control_port_translator:uav_read
	wire  [31:0] spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata;                // SPI_MEDIATOR_spi_control_port_translator:uav_readdata -> SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // SPI_MEDIATOR_spi_control_port_translator:uav_readdatavalid -> SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SPI_MEDIATOR_spi_control_port_translator:uav_debugaccess
	wire   [3:0] spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable;              // SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:m0_byteenable -> SPI_MEDIATOR_spi_control_port_translator:uav_byteenable
	wire         spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid;            // SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_valid -> SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [85:0] spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data;             // SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_data -> SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready;            // SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [85:0] spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         niosii_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                // NIOSII_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         niosii_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                      // NIOSII_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         niosii_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;              // NIOSII_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [94:0] niosii_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                       // NIOSII_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         niosii_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                      // addr_router:sink_ready -> NIOSII_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         niosii_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                       // NIOSII_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire         niosii_data_master_translator_avalon_universal_master_0_agent_cp_valid;                             // NIOSII_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire         niosii_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                     // NIOSII_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [94:0] niosii_data_master_translator_avalon_universal_master_0_agent_cp_data;                              // NIOSII_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire         niosii_data_master_translator_avalon_universal_master_0_agent_cp_ready;                             // addr_router_001:sink_ready -> NIOSII_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                  // NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                        // NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                // NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [94:0] niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                         // NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                        // id_router:sink_ready -> NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire         bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // BRIDGE_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid;                                       // BRIDGE_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // BRIDGE_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [94:0] bridge_s0_translator_avalon_universal_slave_0_agent_rp_data;                                        // BRIDGE_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_001:sink_ready -> BRIDGE_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire         bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket;                                // BRIDGE_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire         bridge_m0_translator_avalon_universal_master_0_agent_cp_valid;                                      // BRIDGE_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire         bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket;                              // BRIDGE_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire  [84:0] bridge_m0_translator_avalon_universal_master_0_agent_cp_data;                                       // BRIDGE_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire         bridge_m0_translator_avalon_universal_master_0_agent_cp_ready;                                      // addr_router_002:sink_ready -> BRIDGE_m0_translator_avalon_universal_master_0_agent:cp_ready
	wire         onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire         onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                   // ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire         onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [84:0] onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_data;                                    // ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire         onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_002:sink_ready -> ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;               // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                     // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;             // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [84:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                      // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                     // id_router_003:sink_ready -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // TIMER_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire         timer_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // TIMER_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire         timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // TIMER_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [84:0] timer_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // TIMER_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire         timer_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_004:sink_ready -> TIMER_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire         spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid;                   // SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire         spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [84:0] spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data;                    // SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire         spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_005:sink_ready -> SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:rp_ready
	wire         addr_router_002_src_endofpacket;                                                                    // addr_router_002:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire         addr_router_002_src_valid;                                                                          // addr_router_002:src_valid -> limiter:cmd_sink_valid
	wire         addr_router_002_src_startofpacket;                                                                  // addr_router_002:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [84:0] addr_router_002_src_data;                                                                           // addr_router_002:src_data -> limiter:cmd_sink_data
	wire   [3:0] addr_router_002_src_channel;                                                                        // addr_router_002:src_channel -> limiter:cmd_sink_channel
	wire         addr_router_002_src_ready;                                                                          // limiter:cmd_sink_ready -> addr_router_002:src_ready
	wire         limiter_rsp_src_endofpacket;                                                                        // limiter:rsp_src_endofpacket -> BRIDGE_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_rsp_src_valid;                                                                              // limiter:rsp_src_valid -> BRIDGE_m0_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_rsp_src_startofpacket;                                                                      // limiter:rsp_src_startofpacket -> BRIDGE_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [84:0] limiter_rsp_src_data;                                                                               // limiter:rsp_src_data -> BRIDGE_m0_translator_avalon_universal_master_0_agent:rp_data
	wire   [3:0] limiter_rsp_src_channel;                                                                            // limiter:rsp_src_channel -> BRIDGE_m0_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_rsp_src_ready;                                                                              // BRIDGE_m0_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire         rst_controller_reset_out_reset;                                                                     // rst_controller:reset_out -> [BRIDGE:reset, BRIDGE_m0_translator:reset, BRIDGE_m0_translator_avalon_universal_master_0_agent:reset, BRIDGE_s0_translator:reset, BRIDGE_s0_translator_avalon_universal_slave_0_agent:reset, BRIDGE_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, JTAG_UART:rst_n, JTAG_UART_avalon_jtag_slave_translator:reset, JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, NIOSII:reset_n, NIOSII_data_master_translator:reset, NIOSII_data_master_translator_avalon_universal_master_0_agent:reset, NIOSII_instruction_master_translator:reset, NIOSII_instruction_master_translator_avalon_universal_master_0_agent:reset, NIOSII_jtag_debug_module_translator:reset, NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, ONCHIP_RAM:reset, ONCHIP_RAM_s1_translator:reset, ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:reset, ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, SPI_MEDIATOR:reset_n, SPI_MEDIATOR_spi_control_port_translator:reset, SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:reset, SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, TIMER:reset_n, TIMER_s1_translator:reset, TIMER_s1_translator_avalon_universal_slave_0_agent:reset, TIMER_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, addr_router_001:reset, addr_router_002:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_002:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, irq_mapper:reset, limiter:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, rsp_xbar_mux_002:reset]
	wire         rst_controller_reset_out_reset_req;                                                                 // rst_controller:reset_req -> ONCHIP_RAM:reset_req
	wire         cmd_xbar_demux_src0_endofpacket;                                                                    // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                          // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                                  // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_src0_data;                                                                           // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [1:0] cmd_xbar_demux_src0_channel;                                                                        // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire         cmd_xbar_demux_src0_ready;                                                                          // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire         cmd_xbar_demux_src1_endofpacket;                                                                    // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                                          // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                                  // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [94:0] cmd_xbar_demux_src1_data;                                                                           // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire   [1:0] cmd_xbar_demux_src1_channel;                                                                        // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire         cmd_xbar_demux_src1_ready;                                                                          // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire         cmd_xbar_demux_001_src0_endofpacket;                                                                // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire         cmd_xbar_demux_001_src0_valid;                                                                      // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire         cmd_xbar_demux_001_src0_startofpacket;                                                              // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_001_src0_data;                                                                       // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [1:0] cmd_xbar_demux_001_src0_channel;                                                                    // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire         cmd_xbar_demux_001_src0_ready;                                                                      // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire         cmd_xbar_demux_001_src1_endofpacket;                                                                // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire         cmd_xbar_demux_001_src1_valid;                                                                      // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire         cmd_xbar_demux_001_src1_startofpacket;                                                              // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [94:0] cmd_xbar_demux_001_src1_data;                                                                       // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire   [1:0] cmd_xbar_demux_001_src1_channel;                                                                    // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire         cmd_xbar_demux_001_src1_ready;                                                                      // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire         rsp_xbar_demux_src0_endofpacket;                                                                    // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                          // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                                  // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [94:0] rsp_xbar_demux_src0_data;                                                                           // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [1:0] rsp_xbar_demux_src0_channel;                                                                        // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                                          // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_src1_endofpacket;                                                                    // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire         rsp_xbar_demux_src1_valid;                                                                          // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire         rsp_xbar_demux_src1_startofpacket;                                                                  // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [94:0] rsp_xbar_demux_src1_data;                                                                           // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire   [1:0] rsp_xbar_demux_src1_channel;                                                                        // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire         rsp_xbar_demux_src1_ready;                                                                          // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                                // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                                      // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                              // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [94:0] rsp_xbar_demux_001_src0_data;                                                                       // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [1:0] rsp_xbar_demux_001_src0_channel;                                                                    // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                                      // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_001_src1_endofpacket;                                                                // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire         rsp_xbar_demux_001_src1_valid;                                                                      // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire         rsp_xbar_demux_001_src1_startofpacket;                                                              // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [94:0] rsp_xbar_demux_001_src1_data;                                                                       // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire   [1:0] rsp_xbar_demux_001_src1_channel;                                                                    // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire         rsp_xbar_demux_001_src1_ready;                                                                      // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire         addr_router_src_endofpacket;                                                                        // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         addr_router_src_valid;                                                                              // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire         addr_router_src_startofpacket;                                                                      // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [94:0] addr_router_src_data;                                                                               // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire   [1:0] addr_router_src_channel;                                                                            // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire         addr_router_src_ready;                                                                              // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                                       // rsp_xbar_mux:src_endofpacket -> NIOSII_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                             // rsp_xbar_mux:src_valid -> NIOSII_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                                     // rsp_xbar_mux:src_startofpacket -> NIOSII_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [94:0] rsp_xbar_mux_src_data;                                                                              // rsp_xbar_mux:src_data -> NIOSII_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [1:0] rsp_xbar_mux_src_channel;                                                                           // rsp_xbar_mux:src_channel -> NIOSII_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_src_ready;                                                                             // NIOSII_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	wire         addr_router_001_src_endofpacket;                                                                    // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire         addr_router_001_src_valid;                                                                          // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire         addr_router_001_src_startofpacket;                                                                  // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [94:0] addr_router_001_src_data;                                                                           // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire   [1:0] addr_router_001_src_channel;                                                                        // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire         addr_router_001_src_ready;                                                                          // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire         rsp_xbar_mux_001_src_endofpacket;                                                                   // rsp_xbar_mux_001:src_endofpacket -> NIOSII_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_001_src_valid;                                                                         // rsp_xbar_mux_001:src_valid -> NIOSII_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_001_src_startofpacket;                                                                 // rsp_xbar_mux_001:src_startofpacket -> NIOSII_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [94:0] rsp_xbar_mux_001_src_data;                                                                          // rsp_xbar_mux_001:src_data -> NIOSII_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [1:0] rsp_xbar_mux_001_src_channel;                                                                       // rsp_xbar_mux_001:src_channel -> NIOSII_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_001_src_ready;                                                                         // NIOSII_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire         cmd_xbar_mux_src_endofpacket;                                                                       // cmd_xbar_mux:src_endofpacket -> NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_src_valid;                                                                             // cmd_xbar_mux:src_valid -> NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_src_startofpacket;                                                                     // cmd_xbar_mux:src_startofpacket -> NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_src_data;                                                                              // cmd_xbar_mux:src_data -> NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [1:0] cmd_xbar_mux_src_channel;                                                                           // cmd_xbar_mux:src_channel -> NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_src_ready;                                                                             // NIOSII_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire         id_router_src_endofpacket;                                                                          // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                                // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                        // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [94:0] id_router_src_data;                                                                                 // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [1:0] id_router_src_channel;                                                                              // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                                // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_mux_001_src_endofpacket;                                                                   // cmd_xbar_mux_001:src_endofpacket -> BRIDGE_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_001_src_valid;                                                                         // cmd_xbar_mux_001:src_valid -> BRIDGE_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_001_src_startofpacket;                                                                 // cmd_xbar_mux_001:src_startofpacket -> BRIDGE_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [94:0] cmd_xbar_mux_001_src_data;                                                                          // cmd_xbar_mux_001:src_data -> BRIDGE_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [1:0] cmd_xbar_mux_001_src_channel;                                                                       // cmd_xbar_mux_001:src_channel -> BRIDGE_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_001_src_ready;                                                                         // BRIDGE_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire         id_router_001_src_endofpacket;                                                                      // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         id_router_001_src_valid;                                                                            // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire         id_router_001_src_startofpacket;                                                                    // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [94:0] id_router_001_src_data;                                                                             // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [1:0] id_router_001_src_channel;                                                                          // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire         id_router_001_src_ready;                                                                            // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire         cmd_xbar_demux_002_src0_endofpacket;                                                                // cmd_xbar_demux_002:src0_endofpacket -> ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_002_src0_valid;                                                                      // cmd_xbar_demux_002:src0_valid -> ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_002_src0_startofpacket;                                                              // cmd_xbar_demux_002:src0_startofpacket -> ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [84:0] cmd_xbar_demux_002_src0_data;                                                                       // cmd_xbar_demux_002:src0_data -> ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [3:0] cmd_xbar_demux_002_src0_channel;                                                                    // cmd_xbar_demux_002:src0_channel -> ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_002_src1_endofpacket;                                                                // cmd_xbar_demux_002:src1_endofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_002_src1_valid;                                                                      // cmd_xbar_demux_002:src1_valid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_002_src1_startofpacket;                                                              // cmd_xbar_demux_002:src1_startofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [84:0] cmd_xbar_demux_002_src1_data;                                                                       // cmd_xbar_demux_002:src1_data -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [3:0] cmd_xbar_demux_002_src1_channel;                                                                    // cmd_xbar_demux_002:src1_channel -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_002_src2_endofpacket;                                                                // cmd_xbar_demux_002:src2_endofpacket -> TIMER_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_002_src2_valid;                                                                      // cmd_xbar_demux_002:src2_valid -> TIMER_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_002_src2_startofpacket;                                                              // cmd_xbar_demux_002:src2_startofpacket -> TIMER_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [84:0] cmd_xbar_demux_002_src2_data;                                                                       // cmd_xbar_demux_002:src2_data -> TIMER_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [3:0] cmd_xbar_demux_002_src2_channel;                                                                    // cmd_xbar_demux_002:src2_channel -> TIMER_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_002_src3_endofpacket;                                                                // cmd_xbar_demux_002:src3_endofpacket -> SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_002_src3_valid;                                                                      // cmd_xbar_demux_002:src3_valid -> SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_002_src3_startofpacket;                                                              // cmd_xbar_demux_002:src3_startofpacket -> SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [84:0] cmd_xbar_demux_002_src3_data;                                                                       // cmd_xbar_demux_002:src3_data -> SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:cp_data
	wire   [3:0] cmd_xbar_demux_002_src3_channel;                                                                    // cmd_xbar_demux_002:src3_channel -> SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rsp_xbar_demux_002_src0_endofpacket;                                                                // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux_002:sink0_endofpacket
	wire         rsp_xbar_demux_002_src0_valid;                                                                      // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux_002:sink0_valid
	wire         rsp_xbar_demux_002_src0_startofpacket;                                                              // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux_002:sink0_startofpacket
	wire  [84:0] rsp_xbar_demux_002_src0_data;                                                                       // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux_002:sink0_data
	wire   [3:0] rsp_xbar_demux_002_src0_channel;                                                                    // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux_002:sink0_channel
	wire         rsp_xbar_demux_002_src0_ready;                                                                      // rsp_xbar_mux_002:sink0_ready -> rsp_xbar_demux_002:src0_ready
	wire         rsp_xbar_demux_003_src0_endofpacket;                                                                // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_002:sink1_endofpacket
	wire         rsp_xbar_demux_003_src0_valid;                                                                      // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_002:sink1_valid
	wire         rsp_xbar_demux_003_src0_startofpacket;                                                              // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_002:sink1_startofpacket
	wire  [84:0] rsp_xbar_demux_003_src0_data;                                                                       // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_002:sink1_data
	wire   [3:0] rsp_xbar_demux_003_src0_channel;                                                                    // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_002:sink1_channel
	wire         rsp_xbar_demux_003_src0_ready;                                                                      // rsp_xbar_mux_002:sink1_ready -> rsp_xbar_demux_003:src0_ready
	wire         rsp_xbar_demux_004_src0_endofpacket;                                                                // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_002:sink2_endofpacket
	wire         rsp_xbar_demux_004_src0_valid;                                                                      // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_002:sink2_valid
	wire         rsp_xbar_demux_004_src0_startofpacket;                                                              // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_002:sink2_startofpacket
	wire  [84:0] rsp_xbar_demux_004_src0_data;                                                                       // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_002:sink2_data
	wire   [3:0] rsp_xbar_demux_004_src0_channel;                                                                    // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_002:sink2_channel
	wire         rsp_xbar_demux_004_src0_ready;                                                                      // rsp_xbar_mux_002:sink2_ready -> rsp_xbar_demux_004:src0_ready
	wire         rsp_xbar_demux_005_src0_endofpacket;                                                                // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_002:sink3_endofpacket
	wire         rsp_xbar_demux_005_src0_valid;                                                                      // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_002:sink3_valid
	wire         rsp_xbar_demux_005_src0_startofpacket;                                                              // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_002:sink3_startofpacket
	wire  [84:0] rsp_xbar_demux_005_src0_data;                                                                       // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_002:sink3_data
	wire   [3:0] rsp_xbar_demux_005_src0_channel;                                                                    // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_002:sink3_channel
	wire         rsp_xbar_demux_005_src0_ready;                                                                      // rsp_xbar_mux_002:sink3_ready -> rsp_xbar_demux_005:src0_ready
	wire         limiter_cmd_src_endofpacket;                                                                        // limiter:cmd_src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire         limiter_cmd_src_startofpacket;                                                                      // limiter:cmd_src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire  [84:0] limiter_cmd_src_data;                                                                               // limiter:cmd_src_data -> cmd_xbar_demux_002:sink_data
	wire   [3:0] limiter_cmd_src_channel;                                                                            // limiter:cmd_src_channel -> cmd_xbar_demux_002:sink_channel
	wire         limiter_cmd_src_ready;                                                                              // cmd_xbar_demux_002:sink_ready -> limiter:cmd_src_ready
	wire         rsp_xbar_mux_002_src_endofpacket;                                                                   // rsp_xbar_mux_002:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire         rsp_xbar_mux_002_src_valid;                                                                         // rsp_xbar_mux_002:src_valid -> limiter:rsp_sink_valid
	wire         rsp_xbar_mux_002_src_startofpacket;                                                                 // rsp_xbar_mux_002:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [84:0] rsp_xbar_mux_002_src_data;                                                                          // rsp_xbar_mux_002:src_data -> limiter:rsp_sink_data
	wire   [3:0] rsp_xbar_mux_002_src_channel;                                                                       // rsp_xbar_mux_002:src_channel -> limiter:rsp_sink_channel
	wire         rsp_xbar_mux_002_src_ready;                                                                         // limiter:rsp_sink_ready -> rsp_xbar_mux_002:src_ready
	wire         cmd_xbar_demux_002_src0_ready;                                                                      // ONCHIP_RAM_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src0_ready
	wire         id_router_002_src_endofpacket;                                                                      // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire         id_router_002_src_valid;                                                                            // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire         id_router_002_src_startofpacket;                                                                    // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [84:0] id_router_002_src_data;                                                                             // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [3:0] id_router_002_src_channel;                                                                          // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire         id_router_002_src_ready;                                                                            // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire         cmd_xbar_demux_002_src1_ready;                                                                      // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src1_ready
	wire         id_router_003_src_endofpacket;                                                                      // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire         id_router_003_src_valid;                                                                            // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire         id_router_003_src_startofpacket;                                                                    // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [84:0] id_router_003_src_data;                                                                             // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [3:0] id_router_003_src_channel;                                                                          // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire         id_router_003_src_ready;                                                                            // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire         cmd_xbar_demux_002_src2_ready;                                                                      // TIMER_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src2_ready
	wire         id_router_004_src_endofpacket;                                                                      // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire         id_router_004_src_valid;                                                                            // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire         id_router_004_src_startofpacket;                                                                    // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [84:0] id_router_004_src_data;                                                                             // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [3:0] id_router_004_src_channel;                                                                          // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire         id_router_004_src_ready;                                                                            // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire         cmd_xbar_demux_002_src3_ready;                                                                      // SPI_MEDIATOR_spi_control_port_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src3_ready
	wire         id_router_005_src_endofpacket;                                                                      // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire         id_router_005_src_valid;                                                                            // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire         id_router_005_src_startofpacket;                                                                    // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [84:0] id_router_005_src_data;                                                                             // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [3:0] id_router_005_src_channel;                                                                          // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire         id_router_005_src_ready;                                                                            // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire   [3:0] limiter_cmd_valid_data;                                                                             // limiter:cmd_src_valid -> cmd_xbar_demux_002:sink_valid
	wire         irq_mapper_receiver0_irq;                                                                           // JTAG_UART:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                                           // TIMER:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                                           // SPI_MEDIATOR:irq -> irq_mapper:receiver2_irq
	wire  [31:0] niosii_d_irq_irq;                                                                                   // irq_mapper:sender_irq -> NIOSII:d_irq

	nios_flash_interface_NIOSII niosii (
		.clk                                   (clock_50_clk),                                                        //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                     //                   reset_n.reset_n
		.d_address                             (niosii_data_master_address),                                          //               data_master.address
		.d_byteenable                          (niosii_data_master_byteenable),                                       //                          .byteenable
		.d_read                                (niosii_data_master_read),                                             //                          .read
		.d_readdata                            (niosii_data_master_readdata),                                         //                          .readdata
		.d_waitrequest                         (niosii_data_master_waitrequest),                                      //                          .waitrequest
		.d_write                               (niosii_data_master_write),                                            //                          .write
		.d_writedata                           (niosii_data_master_writedata),                                        //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (niosii_data_master_debugaccess),                                      //                          .debugaccess
		.i_address                             (niosii_instruction_master_address),                                   //        instruction_master.address
		.i_read                                (niosii_instruction_master_read),                                      //                          .read
		.i_readdata                            (niosii_instruction_master_readdata),                                  //                          .readdata
		.i_waitrequest                         (niosii_instruction_master_waitrequest),                               //                          .waitrequest
		.d_irq                                 (niosii_d_irq_irq),                                                    //                     d_irq.irq
		.jtag_debug_module_resetrequest        (),                                                                    //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (niosii_jtag_debug_module_translator_avalon_anti_slave_0_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (niosii_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (niosii_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (niosii_jtag_debug_module_translator_avalon_anti_slave_0_read),        //                          .read
		.jtag_debug_module_readdata            (niosii_jtag_debug_module_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (niosii_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (niosii_jtag_debug_module_translator_avalon_anti_slave_0_write),       //                          .write
		.jtag_debug_module_writedata           (niosii_jtag_debug_module_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                                     // custom_instruction_master.readra
	);

	nios_flash_interface_ONCHIP_RAM onchip_ram (
		.clk        (clock_50_clk),                                            //   clk1.clk
		.address    (onchip_ram_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.clken      (onchip_ram_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.chipselect (onchip_ram_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.write      (onchip_ram_s1_translator_avalon_anti_slave_0_write),      //       .write
		.readdata   (onchip_ram_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.writedata  (onchip_ram_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (onchip_ram_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                          // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                       //       .reset_req
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (16),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) bridge (
		.clk              (clock_50_clk),                                           //   clk.clk
		.reset            (rst_controller_reset_out_reset),                         // reset.reset
		.s0_waitrequest   (bridge_s0_translator_avalon_anti_slave_0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (bridge_s0_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.s0_readdatavalid (bridge_s0_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (bridge_s0_translator_avalon_anti_slave_0_burstcount),    //      .burstcount
		.s0_writedata     (bridge_s0_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.s0_address       (bridge_s0_translator_avalon_anti_slave_0_address),       //      .address
		.s0_write         (bridge_s0_translator_avalon_anti_slave_0_write),         //      .write
		.s0_read          (bridge_s0_translator_avalon_anti_slave_0_read),          //      .read
		.s0_byteenable    (bridge_s0_translator_avalon_anti_slave_0_byteenable),    //      .byteenable
		.s0_debugaccess   (bridge_s0_translator_avalon_anti_slave_0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (bridge_m0_waitrequest),                                  //    m0.waitrequest
		.m0_readdata      (bridge_m0_readdata),                                     //      .readdata
		.m0_readdatavalid (bridge_m0_readdatavalid),                                //      .readdatavalid
		.m0_burstcount    (bridge_m0_burstcount),                                   //      .burstcount
		.m0_writedata     (bridge_m0_writedata),                                    //      .writedata
		.m0_address       (bridge_m0_address),                                      //      .address
		.m0_write         (bridge_m0_write),                                        //      .write
		.m0_read          (bridge_m0_read),                                         //      .read
		.m0_byteenable    (bridge_m0_byteenable),                                   //      .byteenable
		.m0_debugaccess   (bridge_m0_debugaccess)                                   //      .debugaccess
	);

	nios_flash_interface_JTAG_UART jtag_uart (
		.clk            (clock_50_clk),                                                           //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                        //             reset.reset_n
		.av_chipselect  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                                //               irq.irq
	);

	nios_flash_interface_TIMER timer (
		.clk        (clock_50_clk),                                       //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    // reset.reset_n
		.address    (timer_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                            //   irq.irq
	);

	nios_flash_interface_SPI_MEDIATOR spi_mediator (
		.clk           (clock_50_clk),                                                            //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                                         //            reset.reset_n
		.data_from_cpu (spi_mediator_spi_control_port_translator_avalon_anti_slave_0_writedata),  // spi_control_port.writedata
		.data_to_cpu   (spi_mediator_spi_control_port_translator_avalon_anti_slave_0_readdata),   //                 .readdata
		.mem_addr      (spi_mediator_spi_control_port_translator_avalon_anti_slave_0_address),    //                 .address
		.read_n        (~spi_mediator_spi_control_port_translator_avalon_anti_slave_0_read),      //                 .read_n
		.spi_select    (spi_mediator_spi_control_port_translator_avalon_anti_slave_0_chipselect), //                 .chipselect
		.write_n       (~spi_mediator_spi_control_port_translator_avalon_anti_slave_0_write),     //                 .write_n
		.irq           (irq_mapper_receiver2_irq),                                                //              irq.irq
		.MISO          (spi_mediator_external_MISO),                                              //         external.export
		.MOSI          (spi_mediator_external_MOSI),                                              //                 .export
		.SCLK          (spi_mediator_external_SCLK),                                              //                 .export
		.SS_n          (spi_mediator_external_SS_n)                                               //                 .export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (26),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (26),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) niosii_instruction_master_translator (
		.clk                      (clock_50_clk),                                                                 //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                               //                     reset.reset
		.uav_address              (niosii_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (niosii_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (niosii_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (niosii_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (niosii_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (niosii_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (niosii_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (niosii_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (niosii_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (niosii_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (niosii_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (niosii_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (niosii_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (niosii_instruction_master_read),                                               //                          .read
		.av_readdata              (niosii_instruction_master_readdata),                                           //                          .readdata
		.av_burstcount            (1'b1),                                                                         //               (terminated)
		.av_byteenable            (4'b1111),                                                                      //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                         //               (terminated)
		.av_begintransfer         (1'b0),                                                                         //               (terminated)
		.av_chipselect            (1'b0),                                                                         //               (terminated)
		.av_readdatavalid         (),                                                                             //               (terminated)
		.av_write                 (1'b0),                                                                         //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                         //               (terminated)
		.av_lock                  (1'b0),                                                                         //               (terminated)
		.av_debugaccess           (1'b0),                                                                         //               (terminated)
		.uav_clken                (),                                                                             //               (terminated)
		.av_clken                 (1'b1),                                                                         //               (terminated)
		.uav_response             (2'b00),                                                                        //               (terminated)
		.av_response              (),                                                                             //               (terminated)
		.uav_writeresponserequest (),                                                                             //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                         //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                         //               (terminated)
		.av_writeresponsevalid    ()                                                                              //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (26),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (26),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (1)
	) niosii_data_master_translator (
		.clk                      (clock_50_clk),                                                          //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                        //                     reset.reset
		.uav_address              (niosii_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (niosii_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (niosii_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (niosii_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (niosii_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (niosii_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (niosii_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (niosii_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (niosii_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (niosii_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (niosii_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (niosii_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (niosii_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (niosii_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (niosii_data_master_read),                                               //                          .read
		.av_readdata              (niosii_data_master_readdata),                                           //                          .readdata
		.av_write                 (niosii_data_master_write),                                              //                          .write
		.av_writedata             (niosii_data_master_writedata),                                          //                          .writedata
		.av_debugaccess           (niosii_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount            (1'b1),                                                                  //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                  //               (terminated)
		.av_begintransfer         (1'b0),                                                                  //               (terminated)
		.av_chipselect            (1'b0),                                                                  //               (terminated)
		.av_readdatavalid         (),                                                                      //               (terminated)
		.av_lock                  (1'b0),                                                                  //               (terminated)
		.uav_clken                (),                                                                      //               (terminated)
		.av_clken                 (1'b1),                                                                  //               (terminated)
		.uav_response             (2'b00),                                                                 //               (terminated)
		.av_response              (),                                                                      //               (terminated)
		.uav_writeresponserequest (),                                                                      //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                  //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                  //               (terminated)
		.av_writeresponsevalid    ()                                                                       //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) niosii_jtag_debug_module_translator (
		.clk                      (clock_50_clk),                                                                        //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                      //                    reset.reset
		.uav_address              (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (niosii_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (niosii_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (niosii_jtag_debug_module_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (niosii_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (niosii_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (niosii_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (niosii_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (niosii_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                                    //              (terminated)
		.av_burstcount            (),                                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                //              (terminated)
		.av_writebyteenable       (),                                                                                    //              (terminated)
		.av_lock                  (),                                                                                    //              (terminated)
		.av_chipselect            (),                                                                                    //              (terminated)
		.av_clken                 (),                                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                                //              (terminated)
		.av_outputenable          (),                                                                                    //              (terminated)
		.uav_response             (),                                                                                    //              (terminated)
		.av_response              (2'b00),                                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (16),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) bridge_s0_translator (
		.clk                      (clock_50_clk),                                                         //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                       //                    reset.reset
		.uav_address              (bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (bridge_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (bridge_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (bridge_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (bridge_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (bridge_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount            (bridge_s0_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable            (bridge_s0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (bridge_s0_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (bridge_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (bridge_s0_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                     //              (terminated)
		.av_beginbursttransfer    (),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                     //              (terminated)
		.av_lock                  (),                                                                     //              (terminated)
		.av_chipselect            (),                                                                     //              (terminated)
		.av_clken                 (),                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                 //              (terminated)
		.av_outputenable          (),                                                                     //              (terminated)
		.uav_response             (),                                                                     //              (terminated)
		.av_response              (2'b00),                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                  //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (16),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (16),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) bridge_m0_translator (
		.clk                      (clock_50_clk),                                                 //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                               //                     reset.reset
		.uav_address              (bridge_m0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (bridge_m0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (bridge_m0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (bridge_m0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (bridge_m0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (bridge_m0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (bridge_m0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (bridge_m0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (bridge_m0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (bridge_m0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (bridge_m0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (bridge_m0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (bridge_m0_waitrequest),                                        //                          .waitrequest
		.av_burstcount            (bridge_m0_burstcount),                                         //                          .burstcount
		.av_byteenable            (bridge_m0_byteenable),                                         //                          .byteenable
		.av_read                  (bridge_m0_read),                                               //                          .read
		.av_readdata              (bridge_m0_readdata),                                           //                          .readdata
		.av_readdatavalid         (bridge_m0_readdatavalid),                                      //                          .readdatavalid
		.av_write                 (bridge_m0_write),                                              //                          .write
		.av_writedata             (bridge_m0_writedata),                                          //                          .writedata
		.av_debugaccess           (bridge_m0_debugaccess),                                        //                          .debugaccess
		.av_beginbursttransfer    (1'b0),                                                         //               (terminated)
		.av_begintransfer         (1'b0),                                                         //               (terminated)
		.av_chipselect            (1'b0),                                                         //               (terminated)
		.av_lock                  (1'b0),                                                         //               (terminated)
		.uav_clken                (),                                                             //               (terminated)
		.av_clken                 (1'b1),                                                         //               (terminated)
		.uav_response             (2'b00),                                                        //               (terminated)
		.av_response              (),                                                             //               (terminated)
		.uav_writeresponserequest (),                                                             //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                         //               (terminated)
		.av_writeresponserequest  (1'b0),                                                         //               (terminated)
		.av_writeresponsevalid    ()                                                              //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_ram_s1_translator (
		.clk                      (clock_50_clk),                                                             //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                           //                    reset.reset
		.uav_address              (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (onchip_ram_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (onchip_ram_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (onchip_ram_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (onchip_ram_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (onchip_ram_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (onchip_ram_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken                 (onchip_ram_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_avalon_jtag_slave_translator (
		.clk                      (clock_50_clk),                                                                           //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                         //                    reset.reset
		.uav_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                                       //              (terminated)
		.av_burstcount            (),                                                                                       //              (terminated)
		.av_byteenable            (),                                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                                       //              (terminated)
		.av_lock                  (),                                                                                       //              (terminated)
		.av_clken                 (),                                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                                   //              (terminated)
		.av_debugaccess           (),                                                                                       //              (terminated)
		.av_outputenable          (),                                                                                       //              (terminated)
		.uav_response             (),                                                                                       //              (terminated)
		.av_response              (2'b00),                                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_s1_translator (
		.clk                      (clock_50_clk),                                                        //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                      //                    reset.reset
		.uav_address              (timer_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (timer_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (timer_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (timer_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (timer_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (timer_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (timer_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                    //              (terminated)
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_byteenable            (),                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) spi_mediator_spi_control_port_translator (
		.clk                      (clock_50_clk),                                                                             //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                           //                    reset.reset
		.uav_address              (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (spi_mediator_spi_control_port_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (spi_mediator_spi_control_port_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (spi_mediator_spi_control_port_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (spi_mediator_spi_control_port_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (spi_mediator_spi_control_port_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (spi_mediator_spi_control_port_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                                         //              (terminated)
		.av_burstcount            (),                                                                                         //              (terminated)
		.av_byteenable            (),                                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                                         //              (terminated)
		.av_lock                  (),                                                                                         //              (terminated)
		.av_clken                 (),                                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                                     //              (terminated)
		.av_debugaccess           (),                                                                                         //              (terminated)
		.av_outputenable          (),                                                                                         //              (terminated)
		.uav_response             (),                                                                                         //              (terminated)
		.av_response              (2'b00),                                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                      //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_BEGIN_BURST           (81),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.PKT_BURST_TYPE_H          (78),
		.PKT_BURST_TYPE_L          (77),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_TRANS_EXCLUSIVE       (67),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (84),
		.PKT_THREAD_ID_H           (85),
		.PKT_THREAD_ID_L           (85),
		.PKT_CACHE_H               (92),
		.PKT_CACHE_L               (89),
		.PKT_DATA_SIDEBAND_H       (80),
		.PKT_DATA_SIDEBAND_L       (80),
		.PKT_QOS_H                 (82),
		.PKT_QOS_L                 (82),
		.PKT_ADDR_SIDEBAND_H       (79),
		.PKT_ADDR_SIDEBAND_L       (79),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.ST_DATA_W                 (95),
		.ST_CHANNEL_W              (2),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) niosii_instruction_master_translator_avalon_universal_master_0_agent (
		.clk                     (clock_50_clk),                                                                          //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.av_address              (niosii_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (niosii_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (niosii_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (niosii_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (niosii_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (niosii_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (niosii_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (niosii_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (niosii_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (niosii_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (niosii_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (niosii_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (niosii_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (niosii_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (niosii_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (niosii_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_src_valid),                                                                //        rp.valid
		.rp_data                 (rsp_xbar_mux_src_data),                                                                 //          .data
		.rp_channel              (rsp_xbar_mux_src_channel),                                                              //          .channel
		.rp_startofpacket        (rsp_xbar_mux_src_startofpacket),                                                        //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_src_endofpacket),                                                          //          .endofpacket
		.rp_ready                (rsp_xbar_mux_src_ready),                                                                //          .ready
		.av_response             (),                                                                                      // (terminated)
		.av_writeresponserequest (1'b0),                                                                                  // (terminated)
		.av_writeresponsevalid   ()                                                                                       // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_BEGIN_BURST           (81),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.PKT_BURST_TYPE_H          (78),
		.PKT_BURST_TYPE_L          (77),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_TRANS_EXCLUSIVE       (67),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (84),
		.PKT_THREAD_ID_H           (85),
		.PKT_THREAD_ID_L           (85),
		.PKT_CACHE_H               (92),
		.PKT_CACHE_L               (89),
		.PKT_DATA_SIDEBAND_H       (80),
		.PKT_DATA_SIDEBAND_L       (80),
		.PKT_QOS_H                 (82),
		.PKT_QOS_L                 (82),
		.PKT_ADDR_SIDEBAND_H       (79),
		.PKT_ADDR_SIDEBAND_L       (79),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.ST_DATA_W                 (95),
		.ST_CHANNEL_W              (2),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) niosii_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (clock_50_clk),                                                                   //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.av_address              (niosii_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (niosii_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (niosii_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (niosii_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (niosii_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (niosii_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (niosii_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (niosii_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (niosii_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (niosii_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (niosii_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (niosii_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (niosii_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (niosii_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (niosii_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (niosii_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_001_src_valid),                                                     //        rp.valid
		.rp_data                 (rsp_xbar_mux_001_src_data),                                                      //          .data
		.rp_channel              (rsp_xbar_mux_001_src_channel),                                                   //          .channel
		.rp_startofpacket        (rsp_xbar_mux_001_src_startofpacket),                                             //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_001_src_endofpacket),                                               //          .endofpacket
		.rp_ready                (rsp_xbar_mux_001_src_ready),                                                     //          .ready
		.av_response             (),                                                                               // (terminated)
		.av_writeresponserequest (1'b0),                                                                           // (terminated)
		.av_writeresponsevalid   ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (84),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (2),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clock_50_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                //       clk_reset.reset
		.m0_address              (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                        //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                        //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                         //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                                //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                  //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                      //                .channel
		.rf_sink_ready           (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clock_50_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                // clk_reset.reset
		.in_data           (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                          // (terminated)
		.csr_readdata      (),                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                          // (terminated)
		.almost_full_data  (),                                                                                              // (terminated)
		.almost_empty_data (),                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                          // (terminated)
		.out_empty         (),                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                          // (terminated)
		.out_error         (),                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                          // (terminated)
		.out_channel       ()                                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (84),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (2),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) bridge_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (clock_50_clk),                                                                   //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                   //                .channel
		.rf_sink_ready           (bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (5),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clock_50_clk),                                                                   //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_BEGIN_BURST           (69),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_TRANS_EXCLUSIVE       (57),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (72),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (73),
		.PKT_THREAD_ID_H           (75),
		.PKT_THREAD_ID_L           (75),
		.PKT_CACHE_H               (82),
		.PKT_CACHE_L               (79),
		.PKT_DATA_SIDEBAND_H       (68),
		.PKT_DATA_SIDEBAND_L       (68),
		.PKT_QOS_H                 (70),
		.PKT_QOS_L                 (70),
		.PKT_ADDR_SIDEBAND_H       (67),
		.PKT_ADDR_SIDEBAND_L       (67),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.ST_DATA_W                 (85),
		.ST_CHANNEL_W              (4),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) bridge_m0_translator_avalon_universal_master_0_agent (
		.clk                     (clock_50_clk),                                                          //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.av_address              (bridge_m0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (bridge_m0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (bridge_m0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (bridge_m0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (bridge_m0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (bridge_m0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (bridge_m0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (bridge_m0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (bridge_m0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (bridge_m0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (bridge_m0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_rsp_src_valid),                                                 //        rp.valid
		.rp_data                 (limiter_rsp_src_data),                                                  //          .data
		.rp_channel              (limiter_rsp_src_channel),                                               //          .channel
		.rp_startofpacket        (limiter_rsp_src_startofpacket),                                         //          .startofpacket
		.rp_endofpacket          (limiter_rsp_src_endofpacket),                                           //          .endofpacket
		.rp_ready                (limiter_rsp_src_ready),                                                 //          .ready
		.av_response             (),                                                                      // (terminated)
		.av_writeresponserequest (1'b0),                                                                  // (terminated)
		.av_writeresponsevalid   ()                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_SRC_ID_H              (72),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (73),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (4),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) onchip_ram_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clock_50_clk),                                                                       //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src0_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src0_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_002_src0_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src0_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src0_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src0_channel),                                                    //                .channel
		.rf_sink_ready           (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clock_50_clk),                                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_SRC_ID_H              (72),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (73),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (4),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clock_50_clk),                                                                                     //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                   //       clk_reset.reset
		.m0_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src1_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src1_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_002_src1_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src1_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src1_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src1_channel),                                                                  //                .channel
		.rf_sink_ready           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clock_50_clk),                                                                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                   // clk_reset.reset
		.in_data           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_SRC_ID_H              (72),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (73),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (4),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) timer_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clock_50_clk),                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (timer_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src2_ready),                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src2_valid),                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_002_src2_data),                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src2_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src2_endofpacket),                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src2_channel),                                               //                .channel
		.rf_sink_ready           (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clock_50_clk),                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.in_data           (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_SRC_ID_H              (72),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (73),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (4),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent (
		.clk                     (clock_50_clk),                                                                                       //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                     //       clk_reset.reset
		.m0_address              (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src3_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src3_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_002_src3_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src3_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src3_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src3_channel),                                                                    //                .channel
		.rf_sink_ready           (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clock_50_clk),                                                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                     // clk_reset.reset
		.in_data           (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	nios_flash_interface_addr_router addr_router (
		.sink_ready         (niosii_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (niosii_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (niosii_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (niosii_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (niosii_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clock_50_clk),                                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                 //       src.ready
		.src_valid          (addr_router_src_valid),                                                                 //          .valid
		.src_data           (addr_router_src_data),                                                                  //          .data
		.src_channel        (addr_router_src_channel),                                                               //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                         //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                            //          .endofpacket
	);

	nios_flash_interface_addr_router addr_router_001 (
		.sink_ready         (niosii_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (niosii_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (niosii_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (niosii_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (niosii_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clock_50_clk),                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                      //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                      //          .valid
		.src_data           (addr_router_001_src_data),                                                       //          .data
		.src_channel        (addr_router_001_src_channel),                                                    //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                 //          .endofpacket
	);

	nios_flash_interface_id_router id_router (
		.sink_ready         (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (niosii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clock_50_clk),                                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                      // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                 //       src.ready
		.src_valid          (id_router_src_valid),                                                                 //          .valid
		.src_data           (id_router_src_data),                                                                  //          .data
		.src_channel        (id_router_src_channel),                                                               //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                         //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                            //          .endofpacket
	);

	nios_flash_interface_id_router id_router_001 (
		.sink_ready         (bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clock_50_clk),                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                              //       src.ready
		.src_valid          (id_router_001_src_valid),                                              //          .valid
		.src_data           (id_router_001_src_data),                                               //          .data
		.src_channel        (id_router_001_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                         //          .endofpacket
	);

	nios_flash_interface_addr_router_002 addr_router_002 (
		.sink_ready         (bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clock_50_clk),                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                             //       src.ready
		.src_valid          (addr_router_002_src_valid),                                             //          .valid
		.src_data           (addr_router_002_src_data),                                              //          .data
		.src_channel        (addr_router_002_src_channel),                                           //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                        //          .endofpacket
	);

	nios_flash_interface_id_router_002 id_router_002 (
		.sink_ready         (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clock_50_clk),                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                  //       src.ready
		.src_valid          (id_router_002_src_valid),                                                  //          .valid
		.src_data           (id_router_002_src_data),                                                   //          .data
		.src_channel        (id_router_002_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                             //          .endofpacket
	);

	nios_flash_interface_id_router_002 id_router_003 (
		.sink_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clock_50_clk),                                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                                //       src.ready
		.src_valid          (id_router_003_src_valid),                                                                //          .valid
		.src_data           (id_router_003_src_data),                                                                 //          .data
		.src_channel        (id_router_003_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                           //          .endofpacket
	);

	nios_flash_interface_id_router_002 id_router_004 (
		.sink_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clock_50_clk),                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                             //       src.ready
		.src_valid          (id_router_004_src_valid),                                             //          .valid
		.src_data           (id_router_004_src_data),                                              //          .data
		.src_channel        (id_router_004_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                        //          .endofpacket
	);

	nios_flash_interface_id_router_002 id_router_005 (
		.sink_ready         (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (spi_mediator_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clock_50_clk),                                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_005_src_valid),                                                                  //          .valid
		.src_data           (id_router_005_src_data),                                                                   //          .data
		.src_channel        (id_router_005_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                             //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (73),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (85),
		.ST_CHANNEL_W              (4),
		.VALID_WIDTH               (4),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (clock_50_clk),                       //       clk.clk
		.reset                  (rst_controller_reset_out_reset),     // clk_reset.reset
		.cmd_sink_ready         (addr_router_002_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_002_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_002_src_data),           //          .data
		.cmd_sink_channel       (addr_router_002_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_002_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_002_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),              //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),               //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),            //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),      //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),        //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_002_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_002_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_002_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_002_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_002_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_002_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),              //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),              //          .valid
		.rsp_src_data           (limiter_rsp_src_data),               //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),            //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),      //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),        //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)              // cmd_valid.data
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (1)
	) rst_controller (
		.reset_in0  (~reset_n_reset_n),                   // reset_in0.reset
		.clk        (clock_50_clk),                       //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req  (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	nios_flash_interface_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clock_50_clk),                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_src_ready),             //      sink.ready
		.sink_channel       (addr_router_src_channel),           //          .channel
		.sink_data          (addr_router_src_data),              //          .data
		.sink_startofpacket (addr_router_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	nios_flash_interface_cmd_xbar_demux cmd_xbar_demux_001 (
		.clk                (clock_50_clk),                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_001_src_ready),             //      sink.ready
		.sink_channel       (addr_router_001_src_channel),           //          .channel
		.sink_data          (addr_router_001_src_data),              //          .data
		.sink_startofpacket (addr_router_001_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_001_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_001_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	nios_flash_interface_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clock_50_clk),                          //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	nios_flash_interface_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (clock_50_clk),                          //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	nios_flash_interface_cmd_xbar_demux rsp_xbar_demux (
		.clk                (clock_50_clk),                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	nios_flash_interface_cmd_xbar_demux rsp_xbar_demux_001 (
		.clk                (clock_50_clk),                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	nios_flash_interface_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clock_50_clk),                          //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	nios_flash_interface_rsp_xbar_mux rsp_xbar_mux_001 (
		.clk                 (clock_50_clk),                          //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	nios_flash_interface_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                (clock_50_clk),                          //        clk.clk
		.reset              (rst_controller_reset_out_reset),        //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),                 //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),               //           .channel
		.sink_data          (limiter_cmd_src_data),                  //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),         //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),           //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),                // sink_valid.data
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_002_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_002_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_002_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_002_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_002_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_002_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_002_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_002_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_002_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_002_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_002_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_002_src2_endofpacket),   //           .endofpacket
		.src3_ready         (cmd_xbar_demux_002_src3_ready),         //       src3.ready
		.src3_valid         (cmd_xbar_demux_002_src3_valid),         //           .valid
		.src3_data          (cmd_xbar_demux_002_src3_data),          //           .data
		.src3_channel       (cmd_xbar_demux_002_src3_channel),       //           .channel
		.src3_startofpacket (cmd_xbar_demux_002_src3_startofpacket), //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_002_src3_endofpacket)    //           .endofpacket
	);

	nios_flash_interface_rsp_xbar_demux_002 rsp_xbar_demux_002 (
		.clk                (clock_50_clk),                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	nios_flash_interface_rsp_xbar_demux_002 rsp_xbar_demux_003 (
		.clk                (clock_50_clk),                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	nios_flash_interface_rsp_xbar_demux_002 rsp_xbar_demux_004 (
		.clk                (clock_50_clk),                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	nios_flash_interface_rsp_xbar_demux_002 rsp_xbar_demux_005 (
		.clk                (clock_50_clk),                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	nios_flash_interface_rsp_xbar_mux_002 rsp_xbar_mux_002 (
		.clk                 (clock_50_clk),                          //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_002_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_002_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_002_src0_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_003_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_004_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_005_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	nios_flash_interface_irq_mapper irq_mapper (
		.clk           (clock_50_clk),                   //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (niosii_d_irq_irq)                //    sender.irq
	);

endmodule
